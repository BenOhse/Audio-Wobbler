--Eingaenge: Start/Stop, Wahlschalter Messdauer
--lineare Rampe und Triger erzeugen, log LUT
--Ausgaenge:log. Rampe, Triggersignal
