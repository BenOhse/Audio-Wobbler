Testbench zu taktgenerator.vhdl
