-- Eingaenge: Sollfrequenz
-- Umrechnung Sollfrequenz-->Phaseninkrement, Phasenakku, Sinus LUT
-- Ausgaenge: Amplitudenwert
