Testbench zu software_pwm.vhdl
