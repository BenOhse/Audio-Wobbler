Testbench zu audio_wobbler.vhdl
