--Testbench zu log_frequenzrampe.vhdl
