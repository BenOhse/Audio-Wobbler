--Eingaenge: Amplitudenwert, (Periodendauer)
--Rampe erzeugen, mit Ampl vergleichen
--Ausgaenge: PWM-Signal
