--50MHz clock rein, 20MHz raus
