--Testbench zu sinusgenerator.vhdl
