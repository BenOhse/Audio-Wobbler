-- Zusammenführen der einzelnen Einheiten und Zuordnung zu Pins
